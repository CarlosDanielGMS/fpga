module tb_ula_8_bits;

logic [7:0] a, b;
logic [3:0] s;
logic m, c_in;

logic [7:0] f;
logic a_eq_b, c_out;
endmodule