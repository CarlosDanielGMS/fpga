module ula_74181
(
    input logic [3:0] a, b, s,
    input logic m, c_in,

    output logic [3:0] f,
    output logic a_eq_b, c_out
);
endmodule